library ieee;
use.std_logic_1164.all;

entity procesador is port (
entradas: in std_logic_vector(9 downto 0);
salidas: out std_logic_vector(9 downto 0
);
